`timescale 1ns/1ps
 
module mux();
 
initial begin
$display("Executed DUT code");
end
 
endmodule